/home/witek/Dokumenty/latex/Sprawozdania/PUC/PUC_567/PUC/mod10.vhd