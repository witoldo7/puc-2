/home/witek/Dokumenty/latex/Sprawozdania/PUC/PUC_567/PUC/decod.vhd