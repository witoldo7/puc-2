library verilog;
use verilog.vl_types.all;
entity cw3_vlg_vec_tst is
end cw3_vlg_vec_tst;
